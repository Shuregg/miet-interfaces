`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 14.11.2023 21:28:33
// Design Name: 
// Module Name: SPI
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

/*
1.	��������� ����������� ����� �������������� ��������� �� ����� ������������� ���������.
2.	����������� ��������� �� ����� Verilog, �������� �������� ������� (I?C/SPI), ��� ������������� IP-core, ��������� ��������� � ������� �������.
3.	��������� �������, ��������� � ��������, - �������� test bench ��� ���������� �������?� ��������� ������ �������� ���������� � ��������� ������ ������� ���������.
 ����������, ����������� � ��������/flash, ����� ���� ������������, �� ������ ��������������� ��������� ��������, ���������� � ����������� ������������.

������� � 2. SPI.
������������ ������: Flash-������ W25Q16, 7-���������� ��-�������, ��������� ������� 74HC595, ������ MPU6000.
������� ��� test bench:
1.	������� 4 ����� ������ �� Flash-������ W25Q16.
2.	������� ���������� ������ �� ������ 7-���������� ������-�����, ������������ ����� ��������� �������� 74HC595.
3.	�������� ������ � Flash-������ W25Q16 �� ������ ������-���� ������.
4.	������� ������ �� Flash-������ W25Q16 �� ������ ������-���� ������, ��������� ������� Fast Read.
5.	������� ���������� ������ �� 7-���������� ����������.
6.	������� ������ �� MPU6000 �� ������� 114-117.
7.	������� ���������� ������ �� 7-���������� ����������.
���������� 7-���������� ���������� �� ���������������� �����, ��������� ���������� - �� ������������ �����.
*/
module SPI(
    input   logic  SCLK_I,
    input   logic  MISO_I,
    
    output  logic  MOSI_O,
    output  logic  SS0_O, //Flash
    output  logic  SS1_O, //8-bit Shift register
    output  logic  SS2_O //sensor
    );
    
    
endmodule
